entity signal_simp is
  Port (
    argA     : in bit;
    argB     : in bit;
    rezultat : out bit
  );

end signal_simp;

architecture Behavioral of signal_simp is

begin


end Behavioral;
