entity signal_simp is
  Port (
    argA     : in  bit_vector(3 downto 0);
    argB     : in  bit_vector(3 downto 0);
    rezultat : out bit_vector(3 downto 0)
  );

end signal_simp;

architecture Behavioral of signal_simp is

begin


end Behavioral;
